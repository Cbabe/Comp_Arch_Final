
`timescale 1ns / 1ps
module Test_SRAM;
 // Inputs
 reg [7:0] dataIn;
 reg [7:0] Addr;
 reg CS;
 reg WE;
 reg RD;
 reg Clk;

 // Outputs
 wire [7:0] dataOut;
endmodule;